module add (input src_reg, input src_reg2, output dest_reg);
    
endmodule